** sch_path: /home/bmott/tt_relative_path_test/xsch/tb/ringOsc/ringOsc_tb.sch
**.subckt ringOsc_tb
x1 net1 GND out ringOsc
* noconn out
V1 net1 GND 1.8
**** begin user architecture code



.control

tran 0.1p 10n

wrdata FILE.csv v(out)

.endc
.saveall


.lib /opt/pdk/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt
**** end user architecture code
**.ends

* expanding   symbol:  ip/ringOsc/ringOsc.sym # of pins=3
** sym_path: /home/bmott/tt_relative_path_test/xsch/ip/ringOsc/ringOsc.sym
** sch_path: /home/bmott/tt_relative_path_test/xsch/ip/ringOsc/ringOsc.sch
.subckt ringOsc VDD VSS out
*.opin out
*.iopin VDD
*.iopin VSS
x1 VDD out net1 VSS inv
x2 VDD net1 net2 VSS inv
x3 VDD net2 out VSS inv
.ends


* expanding   symbol:  ip/inv/inv.sym # of pins=4
** sym_path: /home/bmott/tt_relative_path_test/xsch/ip/inv/inv.sym
** sch_path: /home/bmott/tt_relative_path_test/xsch/ip/inv/inv.sch
.subckt inv VDD in out VSS
*.ipin in
*.opin out
*.iopin VDD
*.iopin VSS
XM2 out in VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0 mult=1
+ m=1
XM11 out in VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0
+ mult=1 m=1
.ends

.GLOBAL GND
.end
